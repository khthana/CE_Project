
--
-- VHDL Program Memory Code 
library ieee;
use ieee.std_logic_1164.all;

entity ROM_1kx14 is
  port ( address : in  std_logic_vector(12 downto 0);
         oe      : in  std_logic;
         dout    : out std_logic_vector(13 downto 0)
       );
end ROM_1kx14;

architecture tb_arm5 of ROM_1kx14 is
subtype adr_range is integer range 0 to 220;
-- declare 1Kx14 ROM
subtype ROM_WORD is std_logic_vector(13 downto 0);
type ROM_TABLE is array (0 to 220) of ROM_WORD;
constant ROM : ROM_TABLE := ROM_TABLE'(
   ROM_WORD'("10100000001001"), -- 00000 2809 
   ROM_WORD'("00000000000000"), -- 00001    0 
   ROM_WORD'("00000000000000"), -- 00002    0 
   ROM_WORD'("00000000000000"), -- 00003    0 
   ROM_WORD'("00000000000000"), -- 00004    0 
   ROM_WORD'("00000000000000"), -- 00005    0 
   ROM_WORD'("00000000000000"), -- 00006    0 
   ROM_WORD'("00000000000000"), -- 00007    0 
   ROM_WORD'("00000000000000"), -- 00008    0 
   ROM_WORD'("01011010000011"), -- 00009 1683 
   ROM_WORD'("11000000000000"), -- 00010 3000 
   ROM_WORD'("00000010000101"), -- 00011   85 
   ROM_WORD'("11000000000000"), -- 00012 3000 
   ROM_WORD'("00000010000110"), -- 00013   86 
   ROM_WORD'("11000000000000"), -- 00014 3000 
   ROM_WORD'("00000010001011"), -- 00015   8b 
   ROM_WORD'("11000000000000"), -- 00016 3000 
   ROM_WORD'("00000010000001"), -- 00017   81 
   ROM_WORD'("01001010000011"), -- 00018 1283 
   ROM_WORD'("11000000000000"), -- 00019 3000 
   ROM_WORD'("00000010000001"), -- 00020   81 
   ROM_WORD'("00000010000101"), -- 00021   85 
   ROM_WORD'("00000010000110"), -- 00022   86 
   ROM_WORD'("11000000000110"), -- 00023 3006 
   ROM_WORD'("00000010000011"), -- 00024   83 
   ROM_WORD'("11000010101111"), -- 00025 30af 
   ROM_WORD'("00000010001111"), -- 00026   8f 
   ROM_WORD'("00110100001111"), -- 00027  d0f 
   ROM_WORD'("00000010001111"), -- 00028   8f 
   ROM_WORD'("00110100001111"), -- 00029  d0f 
   ROM_WORD'("00000010001111"), -- 00030   8f 
   ROM_WORD'("00110100001111"), -- 00031  d0f 
   ROM_WORD'("00000010001111"), -- 00032   8f 
   ROM_WORD'("00110100001111"), -- 00033  d0f 
   ROM_WORD'("00000010001111"), -- 00034   8f 
   ROM_WORD'("00110100001111"), -- 00035  d0f 
   ROM_WORD'("00000010001111"), -- 00036   8f 
   ROM_WORD'("00110100001111"), -- 00037  d0f 
   ROM_WORD'("00000010001111"), -- 00038   8f 
   ROM_WORD'("00110100001111"), -- 00039  d0f 
   ROM_WORD'("00000010001111"), -- 00040   8f 
   ROM_WORD'("00110100001111"), -- 00041  d0f 
   ROM_WORD'("00000010001111"), -- 00042   8f 
   ROM_WORD'("00110100001111"), -- 00043  d0f 
   ROM_WORD'("00000010001111"), -- 00044   8f 
   ROM_WORD'("01100000000011"), -- 00045 1803 
   ROM_WORD'("10100011011000"), -- 00046 28d8 
   ROM_WORD'("01110010000011"), -- 00047 1c83 
   ROM_WORD'("10100011011000"), -- 00048 28d8 
   ROM_WORD'("01110100000011"), -- 00049 1d03 
   ROM_WORD'("10100011011000"), -- 00050 28d8 
   ROM_WORD'("11111001010001"), -- 00051 3e51 
   ROM_WORD'("01110000000011"), -- 00052 1c03 
   ROM_WORD'("10100011011000"), -- 00053 28d8 
   ROM_WORD'("11000000000110"), -- 00054 3006 
   ROM_WORD'("00000010000011"), -- 00055   83 
   ROM_WORD'("11000010101111"), -- 00056 30af 
   ROM_WORD'("00000010001111"), -- 00057   8f 
   ROM_WORD'("00110110001111"), -- 00058  d8f 
   ROM_WORD'("00110110001111"), -- 00059  d8f 
   ROM_WORD'("00110110001111"), -- 00060  d8f 
   ROM_WORD'("00110110001111"), -- 00061  d8f 
   ROM_WORD'("00110110001111"), -- 00062  d8f 
   ROM_WORD'("00110110001111"), -- 00063  d8f 
   ROM_WORD'("00110110001111"), -- 00064  d8f 
   ROM_WORD'("00110110001111"), -- 00065  d8f 
   ROM_WORD'("00110110001111"), -- 00066  d8f 
   ROM_WORD'("01100000000011"), -- 00067 1803 
   ROM_WORD'("10100011011000"), -- 00068 28d8 
   ROM_WORD'("01110010000011"), -- 00069 1c83 
   ROM_WORD'("10100011011000"), -- 00070 28d8 
   ROM_WORD'("01110100000011"), -- 00071 1d03 
   ROM_WORD'("10100011011000"), -- 00072 28d8 
   ROM_WORD'("00100000001111"), -- 00073  80f 
   ROM_WORD'("11111001010001"), -- 00074 3e51 
   ROM_WORD'("01110000000011"), -- 00075 1c03 
   ROM_WORD'("10100011011000"), -- 00076 28d8 
   ROM_WORD'("11000000000110"), -- 00077 3006 
   ROM_WORD'("00000010000011"), -- 00078   83 
   ROM_WORD'("11000000100000"), -- 00079 3020 
   ROM_WORD'("00000010000100"), -- 00080   84 
   ROM_WORD'("11000010101111"), -- 00081 30af 
   ROM_WORD'("00000010000000"), -- 00082   80 
   ROM_WORD'("00110110000000"), -- 00083  d80 
   ROM_WORD'("00110110000000"), -- 00084  d80 
   ROM_WORD'("00110110000000"), -- 00085  d80 
   ROM_WORD'("00110110000000"), -- 00086  d80 
   ROM_WORD'("00110110000000"), -- 00087  d80 
   ROM_WORD'("00110110000000"), -- 00088  d80 
   ROM_WORD'("00110110000000"), -- 00089  d80 
   ROM_WORD'("00110110000000"), -- 00090  d80 
   ROM_WORD'("00110110000000"), -- 00091  d80 
   ROM_WORD'("01100000000011"), -- 00092 1803 
   ROM_WORD'("10100011011000"), -- 00093 28d8 
   ROM_WORD'("01110010000011"), -- 00094 1c83 
   ROM_WORD'("10100011011000"), -- 00095 28d8 
   ROM_WORD'("01110100000011"), -- 00096 1d03 
   ROM_WORD'("10100011011000"), -- 00097 28d8 
   ROM_WORD'("00100000000000"), -- 00098  800 
   ROM_WORD'("11111001010001"), -- 00099 3e51 
   ROM_WORD'("01110000000011"), -- 00100 1c03 
   ROM_WORD'("10100011011000"), -- 00101 28d8 
   ROM_WORD'("11000000000110"), -- 00102 3006 
   ROM_WORD'("00000010000011"), -- 00103   83 
   ROM_WORD'("11000011111010"), -- 00104 30fa 
   ROM_WORD'("00000010001111"), -- 00105   8f 
   ROM_WORD'("00110000001111"), -- 00106  c0f 
   ROM_WORD'("00000010001111"), -- 00107   8f 
   ROM_WORD'("00110000001111"), -- 00108  c0f 
   ROM_WORD'("00000010001111"), -- 00109   8f 
   ROM_WORD'("00110000001111"), -- 00110  c0f 
   ROM_WORD'("00000010001111"), -- 00111   8f 
   ROM_WORD'("00110000001111"), -- 00112  c0f 
   ROM_WORD'("00000010001111"), -- 00113   8f 
   ROM_WORD'("00110000001111"), -- 00114  c0f 
   ROM_WORD'("00000010001111"), -- 00115   8f 
   ROM_WORD'("00110000001111"), -- 00116  c0f 
   ROM_WORD'("00000010001111"), -- 00117   8f 
   ROM_WORD'("00110000001111"), -- 00118  c0f 
   ROM_WORD'("00000010001111"), -- 00119   8f 
   ROM_WORD'("00110000001111"), -- 00120  c0f 
   ROM_WORD'("00000010001111"), -- 00121   8f 
   ROM_WORD'("00110000001111"), -- 00122  c0f 
   ROM_WORD'("00000010001111"), -- 00123   8f 
   ROM_WORD'("01100000000011"), -- 00124 1803 
   ROM_WORD'("10100011011000"), -- 00125 28d8 
   ROM_WORD'("01110010000011"), -- 00126 1c83 
   ROM_WORD'("10100011011000"), -- 00127 28d8 
   ROM_WORD'("01110100000011"), -- 00128 1d03 
   ROM_WORD'("10100011011000"), -- 00129 28d8 
   ROM_WORD'("11111000000110"), -- 00130 3e06 
   ROM_WORD'("01110000000011"), -- 00131 1c03 
   ROM_WORD'("10100011011000"), -- 00132 28d8 
   ROM_WORD'("11000000000110"), -- 00133 3006 
   ROM_WORD'("00000010000011"), -- 00134   83 
   ROM_WORD'("11000011111010"), -- 00135 30fa 
   ROM_WORD'("00000010001111"), -- 00136   8f 
   ROM_WORD'("00110110001111"), -- 00137  d8f 
   ROM_WORD'("00110110001111"), -- 00138  d8f 
   ROM_WORD'("00110110001111"), -- 00139  d8f 
   ROM_WORD'("00110110001111"), -- 00140  d8f 
   ROM_WORD'("00110110001111"), -- 00141  d8f 
   ROM_WORD'("00110110001111"), -- 00142  d8f 
   ROM_WORD'("00110110001111"), -- 00143  d8f 
   ROM_WORD'("00110110001111"), -- 00144  d8f 
   ROM_WORD'("00110110001111"), -- 00145  d8f 
   ROM_WORD'("01100000000011"), -- 00146 1803 
   ROM_WORD'("10100011011000"), -- 00147 28d8 
   ROM_WORD'("01110010000011"), -- 00148 1c83 
   ROM_WORD'("10100011011000"), -- 00149 28d8 
   ROM_WORD'("01110100000011"), -- 00150 1d03 
   ROM_WORD'("10100011011000"), -- 00151 28d8 
   ROM_WORD'("00100000001111"), -- 00152  80f 
   ROM_WORD'("11111000000110"), -- 00153 3e06 
   ROM_WORD'("01110000000011"), -- 00154 1c03 
   ROM_WORD'("10100011011000"), -- 00155 28d8 
   ROM_WORD'("11000000000110"), -- 00156 3006 
   ROM_WORD'("00000010000011"), -- 00157   83 
   ROM_WORD'("11000000100000"), -- 00158 3020 
   ROM_WORD'("00000010000100"), -- 00159   84 
   ROM_WORD'("11000011111010"), -- 00160 30fa 
   ROM_WORD'("00000010000000"), -- 00161   80 
   ROM_WORD'("00110010000000"), -- 00162  c80 
   ROM_WORD'("00110010000000"), -- 00163  c80 
   ROM_WORD'("00110010000000"), -- 00164  c80 
   ROM_WORD'("00110010000000"), -- 00165  c80 
   ROM_WORD'("00110010000000"), -- 00166  c80 
   ROM_WORD'("00110010000000"), -- 00167  c80 
   ROM_WORD'("00110010000000"), -- 00168  c80 
   ROM_WORD'("00110010000000"), -- 00169  c80 
   ROM_WORD'("00110010000000"), -- 00170  c80 
   ROM_WORD'("01100000000011"), -- 00171 1803 
   ROM_WORD'("10100011011000"), -- 00172 28d8 
   ROM_WORD'("01110010000011"), -- 00173 1c83 
   ROM_WORD'("10100011011000"), -- 00174 28d8 
   ROM_WORD'("01110100000011"), -- 00175 1d03 
   ROM_WORD'("10100011011000"), -- 00176 28d8 
   ROM_WORD'("00100000000000"), -- 00177  800 
   ROM_WORD'("11111000000110"), -- 00178 3e06 
   ROM_WORD'("01110000000011"), -- 00179 1c03 
   ROM_WORD'("10100011011000"), -- 00180 28d8 
   ROM_WORD'("11000000000111"), -- 00181 3007 
   ROM_WORD'("00000010000011"), -- 00182   83 
   ROM_WORD'("11000010100101"), -- 00183 30a5 
   ROM_WORD'("00000010001111"), -- 00184   8f 
   ROM_WORD'("00111000001111"), -- 00185  e0f 
   ROM_WORD'("01110000000011"), -- 00186 1c03 
   ROM_WORD'("10100011011000"), -- 00187 28d8 
   ROM_WORD'("01110010000011"), -- 00188 1c83 
   ROM_WORD'("10100011011000"), -- 00189 28d8 
   ROM_WORD'("01110100000011"), -- 00190 1d03 
   ROM_WORD'("10100011011000"), -- 00191 28d8 
   ROM_WORD'("00010000001111"), -- 00192  40f 
   ROM_WORD'("11111000000001"), -- 00193 3e01 
   ROM_WORD'("01110000000011"), -- 00194 1c03 
   ROM_WORD'("10100011011000"), -- 00195 28d8 
   ROM_WORD'("11000000000111"), -- 00196 3007 
   ROM_WORD'("00000010000011"), -- 00197   83 
   ROM_WORD'("11000001011010"), -- 00198 305a 
   ROM_WORD'("00000010001111"), -- 00199   8f 
   ROM_WORD'("00111010001111"), -- 00200  e8f 
   ROM_WORD'("01110000000011"), -- 00201 1c03 
   ROM_WORD'("10100011011000"), -- 00202 28d8 
   ROM_WORD'("01110010000011"), -- 00203 1c83 
   ROM_WORD'("10100011011000"), -- 00204 28d8 
   ROM_WORD'("01110100000011"), -- 00205 1d03 
   ROM_WORD'("10100011011000"), -- 00206 28d8 
   ROM_WORD'("00010000001111"), -- 00207  40f 
   ROM_WORD'("11111000000001"), -- 00208 3e01 
   ROM_WORD'("01110000000011"), -- 00209 1c03 
   ROM_WORD'("10100011011000"), -- 00210 28d8 
   ROM_WORD'("01001010000011"), -- 00211 1283 
   ROM_WORD'("11000011111111"), -- 00212 30ff 
   ROM_WORD'("00000010000101"), -- 00213   85 
   ROM_WORD'("00000010000110"), -- 00214   86 
   ROM_WORD'("10100011010111"), -- 00215 28d7 
   ROM_WORD'("01001010000011"), -- 00216 1283 
   ROM_WORD'("11000011111111"), -- 00217 30ff 
   ROM_WORD'("00000010000101"), -- 00218   85 
   ROM_WORD'("10100011011011"), -- 00219 28db 
   ROM_WORD'("00000000000000")  -- 00220    0 
);


     function to_integer(val : std_logic_vector) return adr_range
     is
             variable sum : adr_range;
             variable tmp : integer range 0 to 8192;
             begin
                     tmp := 1;
                     sum := 0;
                     for i in val'low to val'high loop
                             if val(i) = '1' then
                                     sum := sum +tmp;
                             end if;
                             tmp := tmp + tmp;
                     end loop;
                     return sum;
             end to_integer;

	signal LATCH : std_logic_vector(13 downto 0);
begin
       PROG_MEM:
       process(address)
       begin
            -- Read from the program memory
               LATCH <= ROM(to_integer(address));
       end process;

       CTRL_OUTPUT:
       process(oe)
       begin
               if    oe = '0' then
                       dout <= (others => 'Z');
               else
                      -- Read from the program memory
                       dout <= LATCH;
               end if;
       end process;
end tb_arm5;