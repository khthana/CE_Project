
--
-- VHDL Program Memory Code 
library ieee;
use ieee.std_logic_1164.all;

entity ROM_1kx14 is
  port ( address : in  std_logic_vector(12 downto 0);
         oe      : in  std_logic;
         dout    : out std_logic_vector(13 downto 0)
       );
end ROM_1kx14;

architecture tb_arm1 of ROM_1kx14 is
subtype adr_range is integer range 0 to 151;
-- declare 1Kx14 ROM
subtype ROM_WORD is std_logic_vector(13 downto 0);
type ROM_TABLE is array (0 to 151) of ROM_WORD;
constant ROM : ROM_TABLE := ROM_TABLE'(
   ROM_WORD'("10100000001001"), -- 00000 2809 
   ROM_WORD'("00000000000000"), -- 00001    0 
   ROM_WORD'("00000000000000"), -- 00002    0 
   ROM_WORD'("00000000000000"), -- 00003    0 
   ROM_WORD'("00000000000000"), -- 00004    0 
   ROM_WORD'("00000000000000"), -- 00005    0 
   ROM_WORD'("00000000000000"), -- 00006    0 
   ROM_WORD'("00000000000000"), -- 00007    0 
   ROM_WORD'("00000000000000"), -- 00008    0 
   ROM_WORD'("01011010000011"), -- 00009 1683 
   ROM_WORD'("11000000000000"), -- 00010 3000 
   ROM_WORD'("00000010000101"), -- 00011   85 
   ROM_WORD'("11000000000000"), -- 00012 3000 
   ROM_WORD'("00000010000110"), -- 00013   86 
   ROM_WORD'("11000000000000"), -- 00014 3000 
   ROM_WORD'("00000010001011"), -- 00015   8b 
   ROM_WORD'("11000000000000"), -- 00016 3000
   ROM_WORD'("00000010000001"), -- 00017   81
   ROM_WORD'("01001010000011"), -- 00018 1283 
   ROM_WORD'("11000000000000"), -- 00019 3000 
   ROM_WORD'("00000010000001"), -- 00020   81 
   ROM_WORD'("00000010000101"), -- 00021   85 
   ROM_WORD'("00000010000110"), -- 00022   86 
   ROM_WORD'("11000001111111"), -- 00023 307f 
   ROM_WORD'("00000010001111"), -- 00024   8f 
   ROM_WORD'("11000000000111"), -- 00025 3007 
   ROM_WORD'("00000010000011"), -- 00026   83 
   ROM_WORD'("11000000000000"), -- 00027 3000 
   ROM_WORD'("00011100001111"), -- 00028  70f 
   ROM_WORD'("01100000000011"), -- 00029 1803 
   ROM_WORD'("10100010010011"), -- 00030 2893 
   ROM_WORD'("01100010000011"), -- 00031 1883 
   ROM_WORD'("10100010010011"), -- 00032 2893 
   ROM_WORD'("01100100000011"), -- 00033 1903 
   ROM_WORD'("10100010010011"), -- 00034 2893 
   ROM_WORD'("11111010010000"), -- 00035 3e90 
   ROM_WORD'("01110000000011"), -- 00036 1c03 
   ROM_WORD'("10100010010011"), -- 00037 2893 
   ROM_WORD'("11000001111111"), -- 00038 307f 
   ROM_WORD'("00000010001111"), -- 00039   8f 
   ROM_WORD'("11000000000101"), -- 00040 3005 
   ROM_WORD'("00000010000011"), -- 00041   83 
   ROM_WORD'("11000000001111"), -- 00042 300f 
   ROM_WORD'("00011110001111"), -- 00043  78f 
   ROM_WORD'("01100000000011"), -- 00044 1803 
   ROM_WORD'("10100010010011"), -- 00045 2893 
   ROM_WORD'("01110010000011"), -- 00046 1c83 
   ROM_WORD'("10100010010011"), -- 00047 2893 
   ROM_WORD'("01100100000011"), -- 00048 1903 
   ROM_WORD'("10100010010011"), -- 00049 2893 
   ROM_WORD'("00100000001111"), -- 00050  80f 
   ROM_WORD'("11111010000000"), -- 00051 3e80 
   ROM_WORD'("01110000000011"), -- 00052 1c03 
   ROM_WORD'("10100010010011"), -- 00053 2893 
   ROM_WORD'("11000000000000"), -- 00054 3000 
   ROM_WORD'("00000010001111"), -- 00055   8f 
   ROM_WORD'("11000000000110"), -- 00056 3006 
   ROM_WORD'("00000010000011"), -- 00057   83 
   ROM_WORD'("11000000000000"), -- 00058 3000 
   ROM_WORD'("00011100001111"), -- 00059  70f 
   ROM_WORD'("01100000000011"), -- 00060 1803 
   ROM_WORD'("10100010010011"), -- 00061 2893 
   ROM_WORD'("01100010000011"), -- 00062 1883 
   ROM_WORD'("10100010010011"), -- 00063 2893 
   ROM_WORD'("01110100000011"), -- 00064 1d03 
   ROM_WORD'("10100010010011"), -- 00065 2893 
   ROM_WORD'("11000001111111"), -- 00066 307f 
   ROM_WORD'("00000010001111"), -- 00067   8f 
   ROM_WORD'("11000000000100"), -- 00068 3004 
   ROM_WORD'("00000010000011"), -- 00069   83 
   ROM_WORD'("11000011111111"), -- 00070 30ff 
   ROM_WORD'("00011100001111"), -- 00071  70f 
   ROM_WORD'("01110000000011"), -- 00072 1c03 
   ROM_WORD'("10100010010011"), -- 00073 2893 
   ROM_WORD'("01110010000011"), -- 00074 1c83 
   ROM_WORD'("10100010010011"), -- 00075 2893 
   ROM_WORD'("01100100000011"), -- 00076 1903 
   ROM_WORD'("10100010010011"), -- 00077 2893 
   ROM_WORD'("11000000000111"), -- 00078 3007 
   ROM_WORD'("00000010000011"), -- 00079   83 
   ROM_WORD'("11000000000000"), -- 00080 3000 
   ROM_WORD'("11111011111111"), -- 00081 3eff 
   ROM_WORD'("01100000000011"), -- 00082 1803 
   ROM_WORD'("10100010010011"), -- 00083 2893 
   ROM_WORD'("01100010000011"), -- 00084 1883 
   ROM_WORD'("10100010010011"), -- 00085 2893 
   ROM_WORD'("01100100000011"), -- 00086 1903 
   ROM_WORD'("10100010010011"), -- 00087 2893 
   ROM_WORD'("11000000000100"), -- 00088 3004 
   ROM_WORD'("00000010000011"), -- 00089   83 
   ROM_WORD'("11000011111111"), -- 00090 30ff 
   ROM_WORD'("11111011111111"), -- 00091 3eff 
   ROM_WORD'("01110000000011"), -- 00092 1c03 
   ROM_WORD'("10100010010011"), -- 00093 2893 
   ROM_WORD'("01110010000011"), -- 00094 1c83 
   ROM_WORD'("10100010010011"), -- 00095 2893 
   ROM_WORD'("01100100000011"), -- 00096 1903 
   ROM_WORD'("10100010010011"), -- 00097 2893 
   ROM_WORD'("11000000000111"), -- 00098 3007 
   ROM_WORD'("00000010000011"), -- 00099   83 
   ROM_WORD'("11000000000000"), -- 00100 3000 
   ROM_WORD'("11111000000000"), -- 00101 3e00 
   ROM_WORD'("01100000000011"), -- 00102 1803 
   ROM_WORD'("10100010010011"), -- 00103 2893 
   ROM_WORD'("01100010000011"), -- 00104 1883 
   ROM_WORD'("10100010010011"), -- 00105 2893 
   ROM_WORD'("01110100000011"), -- 00106 1d03 
   ROM_WORD'("10100010010011"), -- 00107 2893 
   ROM_WORD'("11000000000000"), -- 00108 3000 
   ROM_WORD'("00000010000011"), -- 00109   83 
   ROM_WORD'("11000010101010"), -- 00110 30aa 
   ROM_WORD'("11100101010101"), -- 00111 3955 
   ROM_WORD'("01100000000011"), -- 00112 1803 
   ROM_WORD'("10100010010011"), -- 00113 2893 
   ROM_WORD'("01100010000011"), -- 00114 1883 
   ROM_WORD'("10100010010011"), -- 00115 2893 
   ROM_WORD'("01110100000011"), -- 00116 1d03 
   ROM_WORD'("10100010010011"), -- 00117 2893 
   ROM_WORD'("11000000000000"), -- 00118 3000 
   ROM_WORD'("00000010000011"), -- 00119   83 
   ROM_WORD'("11000010101010"), -- 00120 30aa 
   ROM_WORD'("00000010001111"), -- 00121   8f 
   ROM_WORD'("11000001010101"), -- 00122 3055 
   ROM_WORD'("00010100001111"), -- 00123  50f 
   ROM_WORD'("01100000000011"), -- 00124 1803 
   ROM_WORD'("10100010010011"), -- 00125 2893 
   ROM_WORD'("01100010000011"), -- 00126 1883 
   ROM_WORD'("10100010010011"), -- 00127 2893 
   ROM_WORD'("01110100000011"), -- 00128 1d03 
   ROM_WORD'("10100010010011"), -- 00129 2893 
   ROM_WORD'("11000000000000"), -- 00130 3000 
   ROM_WORD'("00000010000011"), -- 00131   83 
   ROM_WORD'("11000010101010"), -- 00132 30aa 
   ROM_WORD'("00000010001111"), -- 00133   8f 
   ROM_WORD'("11000001010101"), -- 00134 3055 
   ROM_WORD'("00010110001111"), -- 00135  58f 
   ROM_WORD'("01100000000011"), -- 00136 1803 
   ROM_WORD'("10100010010011"), -- 00137 2893 
   ROM_WORD'("01100010000011"), -- 00138 1883 
   ROM_WORD'("10100010010011"), -- 00139 2893 
   ROM_WORD'("01110100000011"), -- 00140 1d03 
   ROM_WORD'("10100010010011"), -- 00141 2893 
   ROM_WORD'("01001010000011"), -- 00142 1283 
   ROM_WORD'("11000011111111"), -- 00143 30ff 
   ROM_WORD'("00000010000101"), -- 00144   85 
   ROM_WORD'("00000010000110"), -- 00145   86 
   ROM_WORD'("10100010010010"), -- 00146 2892 
   ROM_WORD'("01001010000011"), -- 00147 1283 
   ROM_WORD'("11000011111111"), -- 00148 30ff 
   ROM_WORD'("00000010000101"), -- 00149   85 
   ROM_WORD'("10100010010110"), -- 00150 2896 
   ROM_WORD'("00000000000000")  -- 00151    0 
);


     function to_integer(val : std_logic_vector) return adr_range
     is
             variable sum : adr_range;
             variable tmp : integer range 0 to 8192;
             begin
                     tmp := 1;
                     sum := 0;
                     for i in val'low to val'high loop
                             if val(i) = '1' then
                                     sum := sum +tmp;
                             end if;
                             tmp := tmp + tmp;
                     end loop;
                     return sum;
             end to_integer;

	signal LATCH : std_logic_vector(13 downto 0);
begin
       PROG_MEM:
       process(address)
       begin
            -- Read from the program memory
               LATCH <= ROM(to_integer(address));
       end process;

       CTRL_OUTPUT:
       process(oe)
       begin
               if    oe = '0' then
                       dout <= (others => 'Z');
               else
                      -- Read from the program memory
                       dout <= LATCH;
               end if;
       end process;
end tb_arm1;
