
--
-- VHDL Program Memory Code 
library ieee;
use ieee.std_logic_1164.all;

entity ROM_1kx14 is
  port ( address : in  std_logic_vector(12 downto 0);
         oe      : in  std_logic;
         dout    : out std_logic_vector(13 downto 0)
       );
end ROM_1kx14;

architecture tb_arm3 of ROM_1kx14 is
subtype adr_range is integer range 0 to 161;
-- declare 1Kx14 ROM
subtype ROM_WORD is std_logic_vector(13 downto 0);
type ROM_TABLE is array (0 to 161) of ROM_WORD;
constant ROM : ROM_TABLE := ROM_TABLE'(
   ROM_WORD'("10100000001001"), -- 00000 2809 
   ROM_WORD'("00000000000000"), -- 00001    0 
   ROM_WORD'("00000000000000"), -- 00002    0 
   ROM_WORD'("00000000000000"), -- 00003    0 
   ROM_WORD'("00000000000000"), -- 00004    0 
   ROM_WORD'("00000000000000"), -- 00005    0 
   ROM_WORD'("00000000000000"), -- 00006    0 
   ROM_WORD'("00000000000000"), -- 00007    0 
   ROM_WORD'("00000000000000"), -- 00008    0 
   ROM_WORD'("01011010000011"), -- 00009 1683 
   ROM_WORD'("11000000000000"), -- 00010 3000 
   ROM_WORD'("00000010000101"), -- 00011   85 
   ROM_WORD'("11000000000000"), -- 00012 3000 
   ROM_WORD'("00000010000110"), -- 00013   86 
   ROM_WORD'("11000000000000"), -- 00014 3000 
   ROM_WORD'("00000010001011"), -- 00015   8b 
   ROM_WORD'("11000000000000"), -- 00016 3000 
   ROM_WORD'("00000010000001"), -- 00017   81 
   ROM_WORD'("01001010000011"), -- 00018 1283 
   ROM_WORD'("11000000000000"), -- 00019 3000 
   ROM_WORD'("00000010000001"), -- 00020   81 
   ROM_WORD'("00000010000101"), -- 00021   85 
   ROM_WORD'("00000010000110"), -- 00022   86 
   ROM_WORD'("11000000000111"), -- 00023 3007 
   ROM_WORD'("00000010000011"), -- 00024   83 
   ROM_WORD'("11000001011010"), -- 00025 305a 
   ROM_WORD'("11101010100101"), -- 00026 3aa5 
   ROM_WORD'("01110000000011"), -- 00027 1c03 
   ROM_WORD'("10100010011101"), -- 00028 289d 
   ROM_WORD'("01110010000011"), -- 00029 1c83 
   ROM_WORD'("10100010011101"), -- 00030 289d 
   ROM_WORD'("01100100000011"), -- 00031 1903 
   ROM_WORD'("10100010011101"), -- 00032 289d 
   ROM_WORD'("11111000000001"), -- 00033 3e01 
   ROM_WORD'("01110000000011"), -- 00034 1c03 
   ROM_WORD'("10100010011101"), -- 00035 289d 
   ROM_WORD'("11000000000000"), -- 00036 3000 
   ROM_WORD'("00000010000011"), -- 00037   83 
   ROM_WORD'("11000000000000"), -- 00038 3000 
   ROM_WORD'("11101000000000"), -- 00039 3a00 
   ROM_WORD'("01100000000011"), -- 00040 1803 
   ROM_WORD'("10100010011101"), -- 00041 289d 
   ROM_WORD'("01100010000011"), -- 00042 1883 
   ROM_WORD'("10100010011101"), -- 00043 289d 
   ROM_WORD'("01110100000011"), -- 00044 1d03 
   ROM_WORD'("10100010011101"), -- 00045 289d 
   ROM_WORD'("11111011111111"), -- 00046 3eff 
   ROM_WORD'("01100000000011"), -- 00047 1803 
   ROM_WORD'("10100010011101"), -- 00048 289d 
   ROM_WORD'("11000000000111"), -- 00049 3007 
   ROM_WORD'("00000010000011"), -- 00050   83 
   ROM_WORD'("11000010100101"), -- 00051 30a5 
   ROM_WORD'("00000010001111"), -- 00052   8f 
   ROM_WORD'("11000001011010"), -- 00053 305a 
   ROM_WORD'("00010000001111"), -- 00054  40f 
   ROM_WORD'("01110000000011"), -- 00055 1c03 
   ROM_WORD'("10100010011101"), -- 00056 289d 
   ROM_WORD'("01110010000011"), -- 00057 1c83 
   ROM_WORD'("10100010011101"), -- 00058 289d 
   ROM_WORD'("01100100000011"), -- 00059 1903 
   ROM_WORD'("10100010011101"), -- 00060 289d 
   ROM_WORD'("11111000000001"), -- 00061 3e01 
   ROM_WORD'("01110000000011"), -- 00062 1c03 
   ROM_WORD'("10100010011101"), -- 00063 289d 
   ROM_WORD'("11000000000111"), -- 00064 3007 
   ROM_WORD'("00000010000011"), -- 00065   83 
   ROM_WORD'("11000001011010"), -- 00066 305a 
   ROM_WORD'("00000010001111"), -- 00067   8f 
   ROM_WORD'("11000010100101"), -- 00068 30a5 
   ROM_WORD'("00010010001111"), -- 00069  48f 
   ROM_WORD'("01110000000011"), -- 00070 1c03 
   ROM_WORD'("10100010011101"), -- 00071 289d 
   ROM_WORD'("01110010000011"), -- 00072 1c83 
   ROM_WORD'("10100010011101"), -- 00073 289d 
   ROM_WORD'("01100100000011"), -- 00074 1903 
   ROM_WORD'("10100010011101"), -- 00075 289d 
   ROM_WORD'("00100000001111"), -- 00076  80f 
   ROM_WORD'("11111000000001"), -- 00077 3e01 
   ROM_WORD'("01110000000011"), -- 00078 1c03 
   ROM_WORD'("10100010011101"), -- 00079 289d 
   ROM_WORD'("11000000000111"), -- 00080 3007 
   ROM_WORD'("00000010000011"), -- 00081   83 
   ROM_WORD'("11000000000000"), -- 00082 3000 
   ROM_WORD'("00000010001111"), -- 00083   8f 
   ROM_WORD'("11000000000000"), -- 00084 3000 
   ROM_WORD'("00010000001111"), -- 00085  40f 
   ROM_WORD'("01110000000011"), -- 00086 1c03 
   ROM_WORD'("10100010011101"), -- 00087 289d 
   ROM_WORD'("01110010000011"), -- 00088 1c83 
   ROM_WORD'("10100010011101"), -- 00089 289d 
   ROM_WORD'("01110100000011"), -- 00090 1d03 
   ROM_WORD'("10100010011101"), -- 00091 289d 
   ROM_WORD'("11111011111111"), -- 00092 3eff 
   ROM_WORD'("01100000000011"), -- 00093 1803 
   ROM_WORD'("10100010011101"), -- 00094 289d 
   ROM_WORD'("11000000000000"), -- 00095 3000 
   ROM_WORD'("00000010000011"), -- 00096   83 
   ROM_WORD'("11000001011010"), -- 00097 305a 
   ROM_WORD'("00000010001111"), -- 00098   8f 
   ROM_WORD'("00000110001111"), -- 00099  18f 
   ROM_WORD'("01100000000011"), -- 00100 1803 
   ROM_WORD'("10100010011101"), -- 00101 289d 
   ROM_WORD'("01100010000011"), -- 00102 1883 
   ROM_WORD'("10100010011101"), -- 00103 289d 
   ROM_WORD'("01110100000011"), -- 00104 1d03 
   ROM_WORD'("10100010011101"), -- 00105 289d 
   ROM_WORD'("00100000001111"), -- 00106  80f 
   ROM_WORD'("11111011111111"), -- 00107 3eff 
   ROM_WORD'("01100000000011"), -- 00108 1803 
   ROM_WORD'("10100010011101"), -- 00109 289d 
   ROM_WORD'("11000000000000"), -- 00110 3000 
   ROM_WORD'("00000010000011"), -- 00111   83 
   ROM_WORD'("11000001011010"), -- 00112 305a 
   ROM_WORD'("00000100000011"), -- 00113  103 
   ROM_WORD'("01100000000011"), -- 00114 1803 
   ROM_WORD'("10100010011101"), -- 00115 289d 
   ROM_WORD'("01100010000011"), -- 00116 1883 
   ROM_WORD'("10100010011101"), -- 00117 289d 
   ROM_WORD'("01110100000011"), -- 00118 1d03 
   ROM_WORD'("10100010011101"), -- 00119 289d 
   ROM_WORD'("11111011111111"), -- 00120 3eff 
   ROM_WORD'("01100000000011"), -- 00121 1803 
   ROM_WORD'("10100010011101"), -- 00122 289d 
   ROM_WORD'("11000000000111"), -- 00123 3007 
   ROM_WORD'("00000010000011"), -- 00124   83 
   ROM_WORD'("11000001011010"), -- 00125 305a 
   ROM_WORD'("00000010001111"), -- 00126   8f 
   ROM_WORD'("00100100001111"), -- 00127  90f 
   ROM_WORD'("01110000000011"), -- 00128 1c03 
   ROM_WORD'("10100010011101"), -- 00129 289d 
   ROM_WORD'("01110010000011"), -- 00130 1c83 
   ROM_WORD'("10100010011101"), -- 00131 289d 
   ROM_WORD'("01100100000011"), -- 00132 1903 
   ROM_WORD'("10100010011101"), -- 00133 289d 
   ROM_WORD'("11111001011011"), -- 00134 3e5b 
   ROM_WORD'("01110100000011"), -- 00135 1d03 
   ROM_WORD'("10100010011101"), -- 00136 289d 
   ROM_WORD'("11000000000000"), -- 00137 3000 
   ROM_WORD'("00000010000011"), -- 00138   83 
   ROM_WORD'("11000011111111"), -- 00139 30ff 
   ROM_WORD'("00000010001111"), -- 00140   8f 
   ROM_WORD'("00100110001111"), -- 00141  98f 
   ROM_WORD'("01100000000011"), -- 00142 1803 
   ROM_WORD'("10100010011101"), -- 00143 289d 
   ROM_WORD'("01100010000011"), -- 00144 1883 
   ROM_WORD'("10100010011101"), -- 00145 289d 
   ROM_WORD'("01110100000011"), -- 00146 1d03 
   ROM_WORD'("10100010011101"), -- 00147 289d 
   ROM_WORD'("00100000001111"), -- 00148  80f 
   ROM_WORD'("11111011111111"), -- 00149 3eff 
   ROM_WORD'("01100000000011"), -- 00150 1803 
   ROM_WORD'("10100010011101"), -- 00151 289d 
   ROM_WORD'("01001010000011"), -- 00152 1283 
   ROM_WORD'("11000011111111"), -- 00153 30ff 
   ROM_WORD'("00000010000101"), -- 00154   85 
   ROM_WORD'("00000010000110"), -- 00155   86 
   ROM_WORD'("10100010011100"), -- 00156 289c 
   ROM_WORD'("01001010000011"), -- 00157 1283 
   ROM_WORD'("11000011111111"), -- 00158 30ff 
   ROM_WORD'("00000010000101"), -- 00159   85 
   ROM_WORD'("10100010100000"), -- 00160 28a0 
   ROM_WORD'("00000000000000")  -- 00161    0 
);


     function to_integer(val : std_logic_vector) return adr_range
     is
             variable sum : adr_range;
             variable tmp : integer range 0 to 8192;
             begin
                     tmp := 1;
                     sum := 0;
                     for i in val'low to val'high loop
                             if val(i) = '1' then
                                     sum := sum +tmp;
                             end if;
                             tmp := tmp + tmp;
                     end loop;
                     return sum;
             end to_integer;

	signal LATCH : std_logic_vector(13 downto 0);
begin
       PROG_MEM:
       process(address)
       begin
            -- Read from the program memory
               LATCH <= ROM(to_integer(address));
       end process;

       CTRL_OUTPUT:
       process(oe)
       begin
               if    oe = '0' then
                       dout <= (others => 'Z');
               else
                      -- Read from the program memory
                       dout <= LATCH;
               end if;
       end process;
end tb_arm3;