
--
-- VHDL Program Memory Code 
library ieee;
use ieee.std_logic_1164.all;

entity ROM_1kx14 is
  port ( address : in  std_logic_vector(12 downto 0);
         oe      : in  std_logic;
         dout    : out std_logic_vector(13 downto 0)
       );
end ROM_1kx14;

architecture tb_bit of ROM_1kx14 is
subtype adr_range is integer range 0 to 184;
-- declare 1Kx14 ROM
subtype ROM_WORD is std_logic_vector(13 downto 0);
type ROM_TABLE is array (0 to 184) of ROM_WORD;
constant ROM : ROM_TABLE := ROM_TABLE'(
   ROM_WORD'("10100000001001"), -- 00000 2809 
   ROM_WORD'("00000000000000"), -- 00001    0 
   ROM_WORD'("00000000000000"), -- 00002    0 
   ROM_WORD'("00000000000000"), -- 00003    0 
   ROM_WORD'("00000000000000"), -- 00004    0 
   ROM_WORD'("00000000000000"), -- 00005    0 
   ROM_WORD'("00000000000000"), -- 00006    0 
   ROM_WORD'("00000000000000"), -- 00007    0 
   ROM_WORD'("00000000000000"), -- 00008    0 
   ROM_WORD'("01011010000011"), -- 00009 1683 
   ROM_WORD'("11000000000000"), -- 00010 3000 
   ROM_WORD'("00000010000101"), -- 00011   85 
   ROM_WORD'("11000000000000"), -- 00012 3000 
   ROM_WORD'("00000010000110"), -- 00013   86 
   ROM_WORD'("11000000000000"), -- 00014 3000 
   ROM_WORD'("00000010001011"), -- 00015   8b 
   ROM_WORD'("11000000000000"), -- 00016 3000 
   ROM_WORD'("00000010000001"), -- 00017   81 
   ROM_WORD'("01001010000011"), -- 00018 1283 
   ROM_WORD'("11000000000000"), -- 00019 3000 
   ROM_WORD'("00000010000001"), -- 00020   81 
   ROM_WORD'("00000010000101"), -- 00021   85 
   ROM_WORD'("00000010000110"), -- 00022   86 
   ROM_WORD'("11000000000111"), -- 00023 3007 
   ROM_WORD'("00000010000011"), -- 00024   83 
   ROM_WORD'("11000011111111"), -- 00025 30ff 
   ROM_WORD'("00000010001111"), -- 00026   8f 
   ROM_WORD'("01000000001111"), -- 00027 100f 
   ROM_WORD'("01110000000011"), -- 00028 1c03 
   ROM_WORD'("10100010110100"), -- 00029 28b4 
   ROM_WORD'("01110010000011"), -- 00030 1c83 
   ROM_WORD'("10100010110100"), -- 00031 28b4 
   ROM_WORD'("01110100000011"), -- 00032 1d03 
   ROM_WORD'("10100010110100"), -- 00033 28b4 
   ROM_WORD'("01100000001111"), -- 00034 180f 
   ROM_WORD'("10100010110100"), -- 00035 28b4 
   ROM_WORD'("01000010001111"), -- 00036 108f 
   ROM_WORD'("01110000000011"), -- 00037 1c03 
   ROM_WORD'("10100010110100"), -- 00038 28b4 
   ROM_WORD'("01110010000011"), -- 00039 1c83 
   ROM_WORD'("10100010110100"), -- 00040 28b4 
   ROM_WORD'("01110100000011"), -- 00041 1d03 
   ROM_WORD'("10100010110100"), -- 00042 28b4 
   ROM_WORD'("01100010001111"), -- 00043 188f 
   ROM_WORD'("10100010110100"), -- 00044 28b4 
   ROM_WORD'("01000100001111"), -- 00045 110f 
   ROM_WORD'("01110000000011"), -- 00046 1c03 
   ROM_WORD'("10100010110100"), -- 00047 28b4 
   ROM_WORD'("01110010000011"), -- 00048 1c83 
   ROM_WORD'("10100010110100"), -- 00049 28b4 
   ROM_WORD'("01110100000011"), -- 00050 1d03 
   ROM_WORD'("10100010110100"), -- 00051 28b4 
   ROM_WORD'("01100100001111"), -- 00052 190f 
   ROM_WORD'("10100010110100"), -- 00053 28b4 
   ROM_WORD'("01000110001111"), -- 00054 118f 
   ROM_WORD'("01110000000011"), -- 00055 1c03 
   ROM_WORD'("10100010110100"), -- 00056 28b4 
   ROM_WORD'("01110010000011"), -- 00057 1c83 
   ROM_WORD'("10100010110100"), -- 00058 28b4 
   ROM_WORD'("01110100000011"), -- 00059 1d03 
   ROM_WORD'("10100010110100"), -- 00060 28b4 
   ROM_WORD'("01100110001111"), -- 00061 198f 
   ROM_WORD'("10100010110100"), -- 00062 28b4 
   ROM_WORD'("01001000001111"), -- 00063 120f 
   ROM_WORD'("01110000000011"), -- 00064 1c03 
   ROM_WORD'("10100010110100"), -- 00065 28b4 
   ROM_WORD'("01110010000011"), -- 00066 1c83 
   ROM_WORD'("10100010110100"), -- 00067 28b4 
   ROM_WORD'("01110100000011"), -- 00068 1d03 
   ROM_WORD'("10100010110100"), -- 00069 28b4 
   ROM_WORD'("01101000001111"), -- 00070 1a0f 
   ROM_WORD'("10100010110100"), -- 00071 28b4 
   ROM_WORD'("01001010001111"), -- 00072 128f 
   ROM_WORD'("01110000000011"), -- 00073 1c03 
   ROM_WORD'("10100010110100"), -- 00074 28b4 
   ROM_WORD'("01110010000011"), -- 00075 1c83 
   ROM_WORD'("10100010110100"), -- 00076 28b4 
   ROM_WORD'("01110100000011"), -- 00077 1d03 
   ROM_WORD'("10100010110100"), -- 00078 28b4 
   ROM_WORD'("01101010001111"), -- 00079 1a8f 
   ROM_WORD'("10100010110100"), -- 00080 28b4 
   ROM_WORD'("01001100001111"), -- 00081 130f 
   ROM_WORD'("01110000000011"), -- 00082 1c03 
   ROM_WORD'("10100010110100"), -- 00083 28b4 
   ROM_WORD'("01110010000011"), -- 00084 1c83 
   ROM_WORD'("10100010110100"), -- 00085 28b4 
   ROM_WORD'("01110100000011"), -- 00086 1d03 
   ROM_WORD'("10100010110100"), -- 00087 28b4 
   ROM_WORD'("01101100001111"), -- 00088 1b0f 
   ROM_WORD'("10100010110100"), -- 00089 28b4 
   ROM_WORD'("01001110001111"), -- 00090 138f 
   ROM_WORD'("01110000000011"), -- 00091 1c03 
   ROM_WORD'("10100010110100"), -- 00092 28b4 
   ROM_WORD'("01110010000011"), -- 00093 1c83 
   ROM_WORD'("10100010110100"), -- 00094 28b4 
   ROM_WORD'("01110100000011"), -- 00095 1d03 
   ROM_WORD'("10100010110100"), -- 00096 28b4 
   ROM_WORD'("01101110001111"), -- 00097 1b8f 
   ROM_WORD'("10100010110100"), -- 00098 28b4 
   ROM_WORD'("11000000000111"), -- 00099 3007 
   ROM_WORD'("00000010000011"), -- 00100   83 
   ROM_WORD'("11000000000000"), -- 00101 3000 
   ROM_WORD'("00000010001111"), -- 00102   8f 
   ROM_WORD'("01010000001111"), -- 00103 140f 
   ROM_WORD'("01110000000011"), -- 00104 1c03 
   ROM_WORD'("10100010110100"), -- 00105 28b4 
   ROM_WORD'("01110010000011"), -- 00106 1c83 
   ROM_WORD'("10100010110100"), -- 00107 28b4 
   ROM_WORD'("01110100000011"), -- 00108 1d03 
   ROM_WORD'("10100010110100"), -- 00109 28b4 
   ROM_WORD'("01110000001111"), -- 00110 1c0f 
   ROM_WORD'("10100010110100"), -- 00111 28b4 
   ROM_WORD'("01010010001111"), -- 00112 148f 
   ROM_WORD'("01110000000011"), -- 00113 1c03 
   ROM_WORD'("10100010110100"), -- 00114 28b4 
   ROM_WORD'("01110010000011"), -- 00115 1c83 
   ROM_WORD'("10100010110100"), -- 00116 28b4 
   ROM_WORD'("01110100000011"), -- 00117 1d03 
   ROM_WORD'("10100010110100"), -- 00118 28b4 
   ROM_WORD'("01110010001111"), -- 00119 1c8f 
   ROM_WORD'("10100010110100"), -- 00120 28b4 
   ROM_WORD'("01010100001111"), -- 00121 150f 
   ROM_WORD'("01110000000011"), -- 00122 1c03 
   ROM_WORD'("10100010110100"), -- 00123 28b4 
   ROM_WORD'("01110010000011"), -- 00124 1c83 
   ROM_WORD'("10100010110100"), -- 00125 28b4 
   ROM_WORD'("01110100000011"), -- 00126 1d03 
   ROM_WORD'("10100010110100"), -- 00127 28b4 
   ROM_WORD'("01110100001111"), -- 00128 1d0f 
   ROM_WORD'("10100010110100"), -- 00129 28b4 
   ROM_WORD'("01010110001111"), -- 00130 158f 
   ROM_WORD'("01110000000011"), -- 00131 1c03 
   ROM_WORD'("10100010110100"), -- 00132 28b4 
   ROM_WORD'("01110010000011"), -- 00133 1c83 
   ROM_WORD'("10100010110100"), -- 00134 28b4 
   ROM_WORD'("01110100000011"), -- 00135 1d03 
   ROM_WORD'("10100010110100"), -- 00136 28b4 
   ROM_WORD'("01110110001111"), -- 00137 1d8f 
   ROM_WORD'("10100010110100"), -- 00138 28b4 
   ROM_WORD'("01011000001111"), -- 00139 160f 
   ROM_WORD'("01110000000011"), -- 00140 1c03 
   ROM_WORD'("10100010110100"), -- 00141 28b4 
   ROM_WORD'("01110010000011"), -- 00142 1c83 
   ROM_WORD'("10100010110100"), -- 00143 28b4 
   ROM_WORD'("01110100000011"), -- 00144 1d03 
   ROM_WORD'("10100010110100"), -- 00145 28b4 
   ROM_WORD'("01111000001111"), -- 00146 1e0f 
   ROM_WORD'("10100010110100"), -- 00147 28b4 
   ROM_WORD'("01011010001111"), -- 00148 168f 
   ROM_WORD'("01110000000011"), -- 00149 1c03 
   ROM_WORD'("10100010110100"), -- 00150 28b4 
   ROM_WORD'("01110010000011"), -- 00151 1c83 
   ROM_WORD'("10100010110100"), -- 00152 28b4 
   ROM_WORD'("01110100000011"), -- 00153 1d03 
   ROM_WORD'("10100010110100"), -- 00154 28b4 
   ROM_WORD'("01111010001111"), -- 00155 1e8f 
   ROM_WORD'("10100010110100"), -- 00156 28b4 
   ROM_WORD'("01011100001111"), -- 00157 170f 
   ROM_WORD'("01110000000011"), -- 00158 1c03 
   ROM_WORD'("10100010110100"), -- 00159 28b4 
   ROM_WORD'("01110010000011"), -- 00160 1c83 
   ROM_WORD'("10100010110100"), -- 00161 28b4 
   ROM_WORD'("01110100000011"), -- 00162 1d03 
   ROM_WORD'("10100010110100"), -- 00163 28b4 
   ROM_WORD'("01111100001111"), -- 00164 1f0f 
   ROM_WORD'("10100010110100"), -- 00165 28b4 
   ROM_WORD'("01011110001111"), -- 00166 178f 
   ROM_WORD'("01110000000011"), -- 00167 1c03 
   ROM_WORD'("10100010110100"), -- 00168 28b4 
   ROM_WORD'("01110010000011"), -- 00169 1c83 
   ROM_WORD'("10100010110100"), -- 00170 28b4 
   ROM_WORD'("01110100000011"), -- 00171 1d03 
   ROM_WORD'("10100010110100"), -- 00172 28b4 
   ROM_WORD'("01111110001111"), -- 00173 1f8f 
   ROM_WORD'("10100010110100"), -- 00174 28b4 
   ROM_WORD'("01001010000011"), -- 00175 1283 
   ROM_WORD'("11000011111111"), -- 00176 30ff 
   ROM_WORD'("00000010000101"), -- 00177   85 
   ROM_WORD'("00000010000110"), -- 00178   86 
   ROM_WORD'("10100010110011"), -- 00179 28b3 
   ROM_WORD'("01001010000011"), -- 00180 1283 
   ROM_WORD'("11000011111111"), -- 00181 30ff 
   ROM_WORD'("00000010000101"), -- 00182   85 
   ROM_WORD'("10100010110111"), -- 00183 28b7 
   ROM_WORD'("00000000000000")  -- 00184    0 
);


     function to_integer(val : std_logic_vector) return adr_range
     is
             variable sum : adr_range;
             variable tmp : integer range 0 to 8192;
             begin
                     tmp := 1;
                     sum := 0;
                     for i in val'low to val'high loop
                             if val(i) = '1' then
                                     sum := sum +tmp;
                             end if;
                             tmp := tmp + tmp;
                     end loop;
                     return sum;
             end to_integer;

	signal LATCH : std_logic_vector(13 downto 0);
begin
       PROG_MEM:
       process(address)
       begin
            -- Read from the program memory
               LATCH <= ROM(to_integer(address));
       end process;

       CTRL_OUTPUT:
       process(oe)
       begin
               if    oe = '0' then
                       dout <= (others => 'Z');
               else
                      -- Read from the program memory
                       dout <= LATCH;
               end if;
       end process;
end tb_bit;