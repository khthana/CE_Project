library ieee;
use ieee.std_logic_1164.all;
library exemplar;
use exemplar.exemplar_1164.all;

entity ROM_64x14 is
  port ( address : in  std_logic_vector(5 downto 0);
         dout    : out std_logic_vector(13 downto 0)
       );
end ROM_64x14;

architecture Test of ROM_64x14 is
-- declare 64x14 ROM
subtype ROM_WORD is std_logic_vector(13 downto 0);
type ROM_TABLE is array (0 to 63) of ROM_WORD;
constant ROM : ROM_TABLE := ROM_TABLE'(
   ROM_WORD'("01011010000011"), -- 00000 1683
   ROM_WORD'("11000000000000"), -- 00001 3000 
   ROM_WORD'("00000010000101"), -- 00002   85 
   ROM_WORD'("11000000000000"), -- 00003 3000 
   ROM_WORD'("00000010000110"), -- 00004   86 
   ROM_WORD'("11000000000000"), -- 00005 3000 
   ROM_WORD'("00000010001011"), -- 00006   8b 
   ROM_WORD'("01001010000011"), -- 00007 1283 
   ROM_WORD'("00000010000101"), -- 00008   85 
   ROM_WORD'("00000010000110"), -- 00009   86 
   ROM_WORD'("00100110000101"), -- 00010  985 
   ROM_WORD'("00100110000110"), -- 00011  986 
   ROM_WORD'("10100000001010"), -- 00012 280a 
   ROM_WORD'("11000011111111"), -- 00013 30ff 
   ROM_WORD'("00000010100001"), -- 00014   a1 
   ROM_WORD'("00101110100001"), -- 00015  ba1 
   ROM_WORD'("10100000001111"), -- 00016 280f 
   ROM_WORD'("00000000001000"), -- 00017    8 
   ROM_WORD'("11000011111111"), -- 00018 30ff 
   ROM_WORD'("00000010100010"), -- 00019   a2 
   ROM_WORD'("00101110100010"), -- 00020  ba2 
   ROM_WORD'("10000000001101"), -- 00021 200d 
   ROM_WORD'("10100000010100"), -- 00022 2814 
   ROM_WORD'("00000000001000"), -- 00023    8 
   ROM_WORD'("11000011111100"), -- 00024 30fc 
   ROM_WORD'("00000010100011"), -- 00025   a3 
   ROM_WORD'("00101110100011"), -- 00026  ba3 
   ROM_WORD'("10000000010010"), -- 00027 2012 
   ROM_WORD'("10100000011010"), -- 00028 281a 
   ROM_WORD'("00000000001000"), -- 00029    8 
   ROM_WORD'("00000000000000"), -- 00030    0 
   ROM_WORD'("00000000000000")  -- 00031    0 
   ROM_WORD'("00000000000000"), -- 00032    0
   ROM_WORD'("00000000000000"), -- 00033    0
   ROM_WORD'("00000000000000"), -- 00034    0
   ROM_WORD'("00000000000000"), -- 00035    0
   ROM_WORD'("00000000000000"), -- 00036    0
   ROM_WORD'("00000000000000"), -- 00037    0
   ROM_WORD'("00000000000000"), -- 00038    0
   ROM_WORD'("00000000000000"), -- 00039    0
   ROM_WORD'("00000000000000"), -- 00040    0
   ROM_WORD'("00000000000000"), -- 00041    0
   ROM_WORD'("00000000000000"), -- 00042    0
   ROM_WORD'("00000000000000"), -- 00043    0
   ROM_WORD'("00000000000000"), -- 00044    0
   ROM_WORD'("00000000000000"), -- 00045    0
   ROM_WORD'("00000000000000"), -- 00046    0
   ROM_WORD'("00000000000000"), -- 00047    0
   ROM_WORD'("00000000000000"), -- 00048    0
   ROM_WORD'("00000000000000"), -- 00049    0
   ROM_WORD'("00000000000000"), -- 00050    0
   ROM_WORD'("00000000000000"), -- 00051    0
   ROM_WORD'("00000000000000"), -- 00052    0
   ROM_WORD'("00000000000000"), -- 00053    0
   ROM_WORD'("00000000000000"), -- 00054    0
   ROM_WORD'("00000000000000"), -- 00055    0
   ROM_WORD'("00000000000000"), -- 00056    0
   ROM_WORD'("00000000000000"), -- 00057    0
   ROM_WORD'("00000000000000"), -- 00058    0
   ROM_WORD'("00000000000000"), -- 00059    0
   ROM_WORD'("00000000000000"), -- 00060    0
   ROM_WORD'("00000000000000"), -- 00061    0
   ROM_WORD'("00000000000000"), -- 00062    0
   ROM_WORD'("00000000000000")  -- 00063    0
);

begin
        -- Read from the program memory
        dout <= ROM(evec2int(address));

end Test;
