
--
-- VHDL Program Memory Code 
library ieee;
use ieee.std_logic_1164.all;

entity ROM_1kx14 is
  port ( address : in  std_logic_vector(12 downto 0);
         oe      : in  std_logic;
         dout    : out std_logic_vector(13 downto 0)
       );
end ROM_1kx14;

architecture tb_b2d of ROM_1kx14 is
subtype adr_range is integer range 0 to 127;
-- declare 1Kx14 ROM
subtype ROM_WORD is std_logic_vector(13 downto 0);
type ROM_TABLE is array (0 to 127) of ROM_WORD;
constant ROM : ROM_TABLE := ROM_TABLE'(
   ROM_WORD'("10100000001001"), -- 00000 2809 
   ROM_WORD'("00000000000000"), -- 00001    0 
   ROM_WORD'("00000000000000"), -- 00002    0 
   ROM_WORD'("00000000000000"), -- 00003    0 
   ROM_WORD'("00000000000000"), -- 00004    0 
   ROM_WORD'("00000000000000"), -- 00005    0 
   ROM_WORD'("00000000000000"), -- 00006    0 
   ROM_WORD'("00000000000000"), -- 00007    0 
   ROM_WORD'("00000000000000"), -- 00008    0 
   ROM_WORD'("01011010000011"), -- 00009 1683 
   ROM_WORD'("11000000000000"), -- 00010 3000 
   ROM_WORD'("00000010000101"), -- 00011   85 
   ROM_WORD'("11000000000000"), -- 00012 3000 
   ROM_WORD'("00000010000110"), -- 00013   86 
   ROM_WORD'("11000000000000"), -- 00014 3000 
   ROM_WORD'("00000010001011"), -- 00015   8b 
   ROM_WORD'("11000000000000"), -- 00016 3000 
   ROM_WORD'("00000010000001"), -- 00017   81 
   ROM_WORD'("01001010000011"), -- 00018 1283 
   ROM_WORD'("11000000000000"), -- 00019 3000 
   ROM_WORD'("00000010000001"), -- 00020   81 
   ROM_WORD'("00000010000101"), -- 00021   85 
   ROM_WORD'("00000010000110"), -- 00022   86 
   ROM_WORD'("11000000000000"), -- 00023 3000 
   ROM_WORD'("00000010010010"), -- 00024   92 
   ROM_WORD'("10000001001110"), -- 00025 204e 
   ROM_WORD'("00100000100001"), -- 00026  821 
   ROM_WORD'("11111011111111"), -- 00027 3eff 
   ROM_WORD'("01100000000011"), -- 00028 1803 
   ROM_WORD'("10100001111011"), -- 00029 287b 
   ROM_WORD'("00100000100010"), -- 00030  822 
   ROM_WORD'("11111011111111"), -- 00031 3eff 
   ROM_WORD'("01100000000011"), -- 00032 1803 
   ROM_WORD'("10100001111011"), -- 00033 287b 
   ROM_WORD'("11000001100100"), -- 00034 3064 
   ROM_WORD'("00000010010010"), -- 00035   92 
   ROM_WORD'("10000001001110"), -- 00036 204e 
   ROM_WORD'("00100000100001"), -- 00037  821 
   ROM_WORD'("11111011111111"), -- 00038 3eff 
   ROM_WORD'("01100000000011"), -- 00039 1803 
   ROM_WORD'("10100001111011"), -- 00040 287b 
   ROM_WORD'("00100000100010"), -- 00041  822 
   ROM_WORD'("11111011111110"), -- 00042 3efe 
   ROM_WORD'("01100000000011"), -- 00043 1803 
   ROM_WORD'("10100001111011"), -- 00044 287b 
   ROM_WORD'("11000011111111"), -- 00045 30ff 
   ROM_WORD'("00000010010010"), -- 00046   92 
   ROM_WORD'("10000001001110"), -- 00047 204e 
   ROM_WORD'("00100000100001"), -- 00048  821 
   ROM_WORD'("11111010101010"), -- 00049 3eaa 
   ROM_WORD'("01100000000011"), -- 00050 1803 
   ROM_WORD'("10100001111011"), -- 00051 287b 
   ROM_WORD'("00100000100010"), -- 00052  822 
   ROM_WORD'("11111011111101"), -- 00053 3efd 
   ROM_WORD'("01100000000011"), -- 00054 1803 
   ROM_WORD'("10100001111011"), -- 00055 287b 
   ROM_WORD'("10100001110110"), -- 00056 2876 
   ROM_WORD'("01011010000011"), -- 00057 1683 
   ROM_WORD'("00100000010110"), -- 00058  816 
   ROM_WORD'("00011100010100"), -- 00059  714 
   ROM_WORD'("00000010001101"), -- 00060   8d 
   ROM_WORD'("11111000000110"), -- 00061 3e06 
   ROM_WORD'("01100010000011"), -- 00062 1883 
   ROM_WORD'("10100001000001"), -- 00063 2841 
   ROM_WORD'("00100000001101"), -- 00064  80d 
   ROM_WORD'("00000010001101"), -- 00065   8d 
   ROM_WORD'("11111001100000"), -- 00066 3e60 
   ROM_WORD'("01100000000011"), -- 00067 1803 
   ROM_WORD'("10100001000110"), -- 00068 2846 
   ROM_WORD'("00100000001101"), -- 00069  80d 
   ROM_WORD'("00000010000000"), -- 00070   80 
   ROM_WORD'("01110000000011"), -- 00071 1c03 
   ROM_WORD'("10100001001101"), -- 00072 284d 
   ROM_WORD'("00101010000100"), -- 00073  a84 
   ROM_WORD'("00101000010101"), -- 00074  a15 
   ROM_WORD'("00000010000000"), -- 00075   80 
   ROM_WORD'("00001110000100"), -- 00076  384 
   ROM_WORD'("00000000001000"), -- 00077    8 
   ROM_WORD'("11000000000000"), -- 00078 3000 
   ROM_WORD'("00000010010000"), -- 00079   90 
   ROM_WORD'("00000010100001"), -- 00080   a1 
   ROM_WORD'("00000010100010"), -- 00081   a2 
   ROM_WORD'("11000000001000"), -- 00082 3008 
   ROM_WORD'("00000010010001"), -- 00083   91 
   ROM_WORD'("00100000010010"), -- 00084  812 
   ROM_WORD'("00000010001110"), -- 00085   8e 
   ROM_WORD'("00110010010010"), -- 00086  c92 
   ROM_WORD'("01110000000011"), -- 00087 1c03 
   ROM_WORD'("10100001100011"), -- 00088 2863 
   ROM_WORD'("00100000100001"), -- 00089  821 
   ROM_WORD'("00000010010100"), -- 00090   94 
   ROM_WORD'("00100000100010"), -- 00091  822 
   ROM_WORD'("00000010010101"), -- 00092   95 
   ROM_WORD'("00100000010000"), -- 00093  810 
   ROM_WORD'("10000001101101"), -- 00094 206d 
   ROM_WORD'("00000010010110"), -- 00095   96 
   ROM_WORD'("11000000100001"), -- 00096 3021 
   ROM_WORD'("00000010000100"), -- 00097   84 
   ROM_WORD'("10000000111001"), -- 00098 2039 
   ROM_WORD'("00101010010000"), -- 00099  a90 
   ROM_WORD'("00101110010001"), -- 00100  b91 
   ROM_WORD'("10100001010110"), -- 00101 2856 
   ROM_WORD'("00100000001110"), -- 00102  80e 
   ROM_WORD'("00000010010010"), -- 00103   92 
   ROM_WORD'("00110110001110"), -- 00104  d8e 
   ROM_WORD'("01110000000011"), -- 00105 1c03 
   ROM_WORD'("10100001101100"), -- 00106 286c 
   ROM_WORD'("00101010100010"), -- 00107  aa2 
   ROM_WORD'("00000000001000"), -- 00108    8 
   ROM_WORD'("00011110000010"), -- 00109  782 
   ROM_WORD'("11010000000001"), -- 00110 3401 
   ROM_WORD'("11010000000010"), -- 00111 3402 
   ROM_WORD'("11010000000100"), -- 00112 3404 
   ROM_WORD'("11010000001000"), -- 00113 3408 
   ROM_WORD'("11010000010110"), -- 00114 3416 
   ROM_WORD'("11010000110010"), -- 00115 3432 
   ROM_WORD'("11010001100100"), -- 00116 3464 
   ROM_WORD'("11010000101000"), -- 00117 3428 
   ROM_WORD'("01001010000011"), -- 00118 1283 
   ROM_WORD'("11000011111111"), -- 00119 30ff 
   ROM_WORD'("00000010000101"), -- 00120   85 
   ROM_WORD'("00000010000110"), -- 00121   86 
   ROM_WORD'("10100001111010"), -- 00122 287a 
   ROM_WORD'("01001010000011"), -- 00123 1283 
   ROM_WORD'("11000011111111"), -- 00124 30ff 
   ROM_WORD'("00000010000101"), -- 00125   85 
   ROM_WORD'("10100001111110"), -- 00126 287e 
   ROM_WORD'("00000000000000")  -- 00127    0 
);


     function to_integer(val : std_logic_vector) return adr_range
     is
             variable sum : adr_range;
             variable tmp : integer range 0 to 8192;
             begin
                     tmp := 1;
                     sum := 0;
                     for i in val'low to val'high loop
                             if val(i) = '1' then
                                     sum := sum +tmp;
                             end if;
                             tmp := tmp + tmp;
                     end loop;
                     return sum;
             end to_integer;

	signal LATCH : std_logic_vector(13 downto 0);
begin
       PROG_MEM:
       process(address)
       begin
            -- Read from the program memory
               LATCH <= ROM(to_integer(address));
       end process;

       CTRL_OUTPUT:
       process(oe)
       begin
               if    oe = '0' then
                       dout <= (others => 'Z');
               else
                      -- Read from the program memory
                       dout <= LATCH;
               end if;
       end process;
end tb_b2d;
