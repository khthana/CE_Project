
--
-- VHDL Program Memory Code 
library ieee;
use ieee.std_logic_1164.all;

entity ROM_1kx14 is
  port ( address : in  std_logic_vector(12 downto 0);
         oe      : in  std_logic;
         dout    : out std_logic_vector(13 downto 0)
       );
end ROM_1kx14;

architecture tb_arm2 of ROM_1kx14 is
subtype adr_range is integer range 0 to 201;
-- declare 1Kx14 ROM
subtype ROM_WORD is std_logic_vector(13 downto 0);
type ROM_TABLE is array (0 to 201) of ROM_WORD;
constant ROM : ROM_TABLE := ROM_TABLE'(
   ROM_WORD'("10100000001001"), -- 00000 2809 
   ROM_WORD'("00000000000000"), -- 00001    0 
   ROM_WORD'("00000000000000"), -- 00002    0 
   ROM_WORD'("00000000000000"), -- 00003    0 
   ROM_WORD'("00000000000000"), -- 00004    0 
   ROM_WORD'("00000000000000"), -- 00005    0 
   ROM_WORD'("00000000000000"), -- 00006    0 
   ROM_WORD'("00000000000000"), -- 00007    0 
   ROM_WORD'("00000000000000"), -- 00008    0 
   ROM_WORD'("01011010000011"), -- 00009 1683 
   ROM_WORD'("11000000000000"), -- 00010 3000 
   ROM_WORD'("00000010000101"), -- 00011   85 
   ROM_WORD'("11000000000000"), -- 00012 3000 
   ROM_WORD'("00000010000110"), -- 00013   86 
   ROM_WORD'("11000000000000"), -- 00014 3000 
   ROM_WORD'("00000010001011"), -- 00015   8b 
   ROM_WORD'("11000000000000"), -- 00016 3000 
   ROM_WORD'("00000010000001"), -- 00017   81 
   ROM_WORD'("01001010000011"), -- 00018 1283 
   ROM_WORD'("11000000000000"), -- 00019 3000 
   ROM_WORD'("00000010000001"), -- 00020   81 
   ROM_WORD'("00000010000101"), -- 00021   85 
   ROM_WORD'("00000010000110"), -- 00022   86 
   ROM_WORD'("11000011111111"), -- 00023 30ff 
   ROM_WORD'("00000010001111"), -- 00024   8f 
   ROM_WORD'("11000000000100"), -- 00025 3004 
   ROM_WORD'("00000010000011"), -- 00026   83 
   ROM_WORD'("11000001111111"), -- 00027 307f 
   ROM_WORD'("00001000001111"), -- 00028  20f 
   ROM_WORD'("01110000000011"), -- 00029 1c03 
   ROM_WORD'("10100011000101"), -- 00030 28c5 
   ROM_WORD'("01110010000011"), -- 00031 1c83 
   ROM_WORD'("10100011000101"), -- 00032 28c5 
   ROM_WORD'("01100100000011"), -- 00033 1903 
   ROM_WORD'("10100011000101"), -- 00034 28c5 
   ROM_WORD'("11111010000000"), -- 00035 3e80 
   ROM_WORD'("01110000000011"), -- 00036 1c03 
   ROM_WORD'("10100011000101"), -- 00037 28c5 
   ROM_WORD'("11000011111111"), -- 00038 30ff 
   ROM_WORD'("00000010001111"), -- 00039   8f 
   ROM_WORD'("11000000000000"), -- 00040 3000 
   ROM_WORD'("00000010000011"), -- 00041   83 
   ROM_WORD'("11000011111111"), -- 00042 30ff 
   ROM_WORD'("00001010001111"), -- 00043  28f 
   ROM_WORD'("01110000000011"), -- 00044 1c03 
   ROM_WORD'("10100011000101"), -- 00045 28c5 
   ROM_WORD'("01110010000011"), -- 00046 1c83 
   ROM_WORD'("10100011000101"), -- 00047 28c5 
   ROM_WORD'("01110100000011"), -- 00048 1d03 
   ROM_WORD'("10100011000101"), -- 00049 28c5 
   ROM_WORD'("11000000000000"), -- 00050 3000 
   ROM_WORD'("00000010001111"), -- 00051   8f 
   ROM_WORD'("11000000000111"), -- 00052 3007 
   ROM_WORD'("00000010000011"), -- 00053   83 
   ROM_WORD'("11000011111111"), -- 00054 30ff 
   ROM_WORD'("00001000001111"), -- 00055  20f 
   ROM_WORD'("01100000000011"), -- 00056 1803 
   ROM_WORD'("10100011000101"), -- 00057 28c5 
   ROM_WORD'("01100010000011"), -- 00058 1883 
   ROM_WORD'("10100011000101"), -- 00059 28c5 
   ROM_WORD'("01100100000011"), -- 00060 1903 
   ROM_WORD'("10100011000101"), -- 00061 28c5 
   ROM_WORD'("11111011111111"), -- 00062 3eff 
   ROM_WORD'("01110000000011"), -- 00063 1c03 
   ROM_WORD'("10100011000101"), -- 00064 28c5 
   ROM_WORD'("11000000000000"), -- 00065 3000 
   ROM_WORD'("00000010001111"), -- 00066   8f 
   ROM_WORD'("11000000000100"), -- 00067 3004 
   ROM_WORD'("00000010000011"), -- 00068   83 
   ROM_WORD'("11000000000001"), -- 00069 3001 
   ROM_WORD'("00001000001111"), -- 00070  20f 
   ROM_WORD'("01100000000011"), -- 00071 1803 
   ROM_WORD'("10100011000101"), -- 00072 28c5 
   ROM_WORD'("01100010000011"), -- 00073 1883 
   ROM_WORD'("10100011000101"), -- 00074 28c5 
   ROM_WORD'("01100100000011"), -- 00075 1903 
   ROM_WORD'("10100011000101"), -- 00076 28c5 
   ROM_WORD'("11111000000001"), -- 00077 3e01 
   ROM_WORD'("01110000000011"), -- 00078 1c03 
   ROM_WORD'("10100011000101"), -- 00079 28c5 
   ROM_WORD'("11000000000100"), -- 00080 3004 
   ROM_WORD'("00000010000011"), -- 00081   83 
   ROM_WORD'("11000001111111"), -- 00082 307f 
   ROM_WORD'("11110011111111"), -- 00083 3cff 
   ROM_WORD'("01110000000011"), -- 00084 1c03 
   ROM_WORD'("10100011000101"), -- 00085 28c5 
   ROM_WORD'("01110010000011"), -- 00086 1c83 
   ROM_WORD'("10100011000101"), -- 00087 28c5 
   ROM_WORD'("01100100000011"), -- 00088 1903 
   ROM_WORD'("10100011000101"), -- 00089 28c5 
   ROM_WORD'("11111010000000"), -- 00090 3e80 
   ROM_WORD'("01110000000011"), -- 00091 1c03 
   ROM_WORD'("10100011000101"), -- 00092 28c5 
   ROM_WORD'("11000000000000"), -- 00093 3000 
   ROM_WORD'("00000010000011"), -- 00094   83 
   ROM_WORD'("11000011111111"), -- 00095 30ff 
   ROM_WORD'("11110011111111"), -- 00096 3cff 
   ROM_WORD'("01110000000011"), -- 00097 1c03 
   ROM_WORD'("10100011000101"), -- 00098 28c5 
   ROM_WORD'("01110010000011"), -- 00099 1c83 
   ROM_WORD'("10100011000101"), -- 00100 28c5 
   ROM_WORD'("01110100000011"), -- 00101 1d03 
   ROM_WORD'("10100011000101"), -- 00102 28c5 
   ROM_WORD'("11000000000111"), -- 00103 3007 
   ROM_WORD'("00000010000011"), -- 00104   83 
   ROM_WORD'("11000011111111"), -- 00105 30ff 
   ROM_WORD'("11110000000000"), -- 00106 3c00 
   ROM_WORD'("01100000000011"), -- 00107 1803 
   ROM_WORD'("10100011000101"), -- 00108 28c5 
   ROM_WORD'("01100010000011"), -- 00109 1883 
   ROM_WORD'("10100011000101"), -- 00110 28c5 
   ROM_WORD'("01100100000011"), -- 00111 1903 
   ROM_WORD'("10100011000101"), -- 00112 28c5 
   ROM_WORD'("11111011111111"), -- 00113 3eff 
   ROM_WORD'("01110000000011"), -- 00114 1c03 
   ROM_WORD'("10100011000101"), -- 00115 28c5 
   ROM_WORD'("11000000000100"), -- 00116 3004 
   ROM_WORD'("00000010000011"), -- 00117   83 
   ROM_WORD'("11000010000001"), -- 00118 3081 
   ROM_WORD'("11110010000000"), -- 00119 3c80 
   ROM_WORD'("01100000000011"), -- 00120 1803 
   ROM_WORD'("10100011000101"), -- 00121 28c5 
   ROM_WORD'("01100010000011"), -- 00122 1883 
   ROM_WORD'("10100011000101"), -- 00123 28c5 
   ROM_WORD'("01100100000011"), -- 00124 1903 
   ROM_WORD'("10100011000101"), -- 00125 28c5 
   ROM_WORD'("11111000000001"), -- 00126 3e01 
   ROM_WORD'("01110000000011"), -- 00127 1c03 
   ROM_WORD'("10100011000101"), -- 00128 28c5 
   ROM_WORD'("11000000000111"), -- 00129 3007 
   ROM_WORD'("00000010000011"), -- 00130   83 
   ROM_WORD'("11000010101010"), -- 00131 30aa 
   ROM_WORD'("11101001010101"), -- 00132 3a55 
   ROM_WORD'("01110000000011"), -- 00133 1c03 
   ROM_WORD'("10100011000101"), -- 00134 28c5 
   ROM_WORD'("01110010000011"), -- 00135 1c83 
   ROM_WORD'("10100011000101"), -- 00136 28c5 
   ROM_WORD'("01100100000011"), -- 00137 1903 
   ROM_WORD'("10100011000101"), -- 00138 28c5 
   ROM_WORD'("11111000000001"), -- 00139 3e01 
   ROM_WORD'("01110000000011"), -- 00140 1c03 
   ROM_WORD'("10100011000101"), -- 00141 28c5 
   ROM_WORD'("11000000000000"), -- 00142 3000 
   ROM_WORD'("00000010000011"), -- 00143   83 
   ROM_WORD'("11000011111111"), -- 00144 30ff 
   ROM_WORD'("11101011111111"), -- 00145 3aff 
   ROM_WORD'("01100000000011"), -- 00146 1803 
   ROM_WORD'("10100011000101"), -- 00147 28c5 
   ROM_WORD'("01100010000011"), -- 00148 1883 
   ROM_WORD'("10100011000101"), -- 00149 28c5 
   ROM_WORD'("01110100000011"), -- 00150 1d03 
   ROM_WORD'("10100011000101"), -- 00151 28c5 
   ROM_WORD'("11000000000111"), -- 00152 3007 
   ROM_WORD'("00000010000011"), -- 00153   83 
   ROM_WORD'("11000001010101"), -- 00154 3055 
   ROM_WORD'("00000010001111"), -- 00155   8f 
   ROM_WORD'("11000010101010"), -- 00156 30aa 
   ROM_WORD'("00011010001111"), -- 00157  68f 
   ROM_WORD'("01110000000011"), -- 00158 1c03 
   ROM_WORD'("10100011000101"), -- 00159 28c5 
   ROM_WORD'("01110010000011"), -- 00160 1c83 
   ROM_WORD'("10100011000101"), -- 00161 28c5 
   ROM_WORD'("01100100000011"), -- 00162 1903 
   ROM_WORD'("10100011000101"), -- 00163 28c5 
   ROM_WORD'("00100000001111"), -- 00164  80f 
   ROM_WORD'("11111000000001"), -- 00165 3e01 
   ROM_WORD'("01110000000011"), -- 00166 1c03 
   ROM_WORD'("10100011000101"), -- 00167 28c5 
   ROM_WORD'("11000000000000"), -- 00168 3000 
   ROM_WORD'("00000010000011"), -- 00169   83 
   ROM_WORD'("11000011111111"), -- 00170 30ff 
   ROM_WORD'("00000010001111"), -- 00171   8f 
   ROM_WORD'("11000011111111"), -- 00172 30ff 
   ROM_WORD'("00011000001111"), -- 00173  60f 
   ROM_WORD'("01100000000011"), -- 00174 1803 
   ROM_WORD'("10100011000101"), -- 00175 28c5 
   ROM_WORD'("01100010000011"), -- 00176 1883 
   ROM_WORD'("10100011000101"), -- 00177 28c5 
   ROM_WORD'("01110100000011"), -- 00178 1d03 
   ROM_WORD'("10100011000101"), -- 00179 28c5 
   ROM_WORD'("11000000000111"), -- 00180 3007 
   ROM_WORD'("00000010000011"), -- 00181   83 
   ROM_WORD'("11000000000000"), -- 00182 3000 
   ROM_WORD'("00000010001111"), -- 00183   8f 
   ROM_WORD'("11000000000000"), -- 00184 3000 
   ROM_WORD'("00011010001111"), -- 00185  68f 
   ROM_WORD'("01110000000011"), -- 00186 1c03 
   ROM_WORD'("10100011000101"), -- 00187 28c5 
   ROM_WORD'("01110010000011"), -- 00188 1c83 
   ROM_WORD'("10100011000101"), -- 00189 28c5 
   ROM_WORD'("01110100000011"), -- 00190 1d03 
   ROM_WORD'("10100011000101"), -- 00191 28c5 
   ROM_WORD'("01001010000011"), -- 00192 1283 
   ROM_WORD'("11000011111111"), -- 00193 30ff 
   ROM_WORD'("00000010000101"), -- 00194   85 
   ROM_WORD'("00000010000110"), -- 00195   86 
   ROM_WORD'("10100011000100"), -- 00196 28c4 
   ROM_WORD'("01001010000011"), -- 00197 1283 
   ROM_WORD'("11000011111111"), -- 00198 30ff 
   ROM_WORD'("00000010000101"), -- 00199   85 
   ROM_WORD'("10100011001000"), -- 00200 28c8 
   ROM_WORD'("00000000000000")  -- 00201    0 
);


     function to_integer(val : std_logic_vector) return adr_range
     is
             variable sum : adr_range;
             variable tmp : integer range 0 to 8192;
             begin
                     tmp := 1;
                     sum := 0;
                     for i in val'low to val'high loop
                             if val(i) = '1' then
                                     sum := sum +tmp;
                             end if;
                             tmp := tmp + tmp;
                     end loop;
                     return sum;
             end to_integer;

	signal LATCH : std_logic_vector(13 downto 0);
begin
       PROG_MEM:
       process(address)
       begin
            -- Read from the program memory
               LATCH <= ROM(to_integer(address));
       end process;

       CTRL_OUTPUT:
       process(oe)
       begin
               if    oe = '0' then
                       dout <= (others => 'Z');
               else
                      -- Read from the program memory
                       dout <= LATCH;
               end if;
       end process;
end tb_arm2;